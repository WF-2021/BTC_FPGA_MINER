//	********************************************************************************
//	ģ������extend_message_calc
//	��  �ܣ�ͨ����Ϣ��M��������չ��Ϣ��W
//	��	Դ��LUT-136��REG-513
//	********************************************************************************
module extend_message_calc # (
	
	//	�������
	parameter		MODULE_INDEX		= 0				,	//	ģ���ţ�0~63
	parameter		WORD_NUM			= 16			,	//	WORD������16
	parameter		DATA_WID			= 32				//	WORDλ��32
	)
	(
	
	//	�����ź�
	input								clk				,	//	ģ�鹤��ʱ���ź�
	input								rst				,	//	clkʱ���򣬸�λ
	input	[WORD_NUM*DATA_WID	-1:0]	iv_m_data		,	//	clkʱ����������Ϣ������M
	input								i_m_data_vld	,	//	clkʱ����������Ϣ������M��Ч
	
	//	����ź�
	output	[WORD_NUM*DATA_WID	-1:0]	ov_m_data		,	//	clkʱ���������Ϣ������M
	output								o_m_data_vld	,	//	clkʱ���������Ϣ������M��Ч
	output	[DATA_WID			-1:0]	ov_w_data		,	//	clkʱ���������չ��Ϣ������W
	output								o_w_data_vld		//	clkʱ���������չ��Ϣ������W��Ч
	);
	
	
	//  ===============================================================================================
	//	�������źš�����˵��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
	//  -----------------------------------------------------------------
	//	rou0����
	//	rou0(x) = s7(x) ^ s18(x) ^ r3(x)
	//  -----------------------------------------------------------------
	function [DATA_WID-1:0] rou0;
		
		//	�����ź�
		input	[DATA_WID	-1:0]	data;
		
		//	�������� 
		reg		[DATA_WID	-1:0]	s7	;
		reg		[DATA_WID	-1:0]	s18	;
		reg		[DATA_WID	-1:0]	r3	;
		
		//	�������  
		begin
			s7		= {data[6:0],	data[DATA_WID-1:7]};
			s18		= {data[17:0],	data[DATA_WID-1:18]};
			r3		= {{(3){1'b0}},	data[DATA_WID-1:3]};
			rou0	= s7 ^ s18 ^ r3;
		end
	endfunction
	
	//  -----------------------------------------------------------------
	//	rou1����
	//	rou1(x) = s17(x) ^ s19(x) ^ r10(x)
	//  -----------------------------------------------------------------
	function [DATA_WID-1:0] rou1;
		
		//	�����ź�
		input	[DATA_WID	-1:0]	data;
		
		//	�������� 
		reg		[DATA_WID	-1:0]	s17;
		reg		[DATA_WID	-1:0]	s19;
		reg		[DATA_WID	-1:0]	r10;
		
		//	�������  
		begin
			s17		= {data[16:0],		data[DATA_WID-1:17]};
			s19		= {data[18:0],		data[DATA_WID-1:19]};
			r10		= {{(10){1'b0}},	data[DATA_WID-1:10]};
			rou1	= s17 ^ s19 ^ r10;
		end
	endfunction
	
	//  -------------------------------------------------------------------------------------
	//	�ź�˵��
	//  -------------------------------------------------------------------------------------
	wire	[DATA_WID	-1:0]	m_data_word		[WORD_NUM	-1:0]	;	//	clkʱ����������Ϣ������M����
	reg		[DATA_WID	-1:0]	m_data_word_reg	[WORD_NUM	-1:0]	;	//	clkʱ������Ϣ������M������
	reg							data_vld_reg	= 1'b0				;	//	clkʱ����������Ϣ������M��Ч����1��

	
	//  ===============================================================================================
	//	��չ��Ϣ��W����
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	������Ϣ������M����
	//	��������Ϣ��M����32bit��wordΪ��λ�����з���
	//  -------------------------------------------------------------------------------------	
	genvar i;	
	generate
		for(i=0; i<WORD_NUM; i=i+1) begin : m_data_word_loop
			assign m_data_word[i] = iv_m_data[(DATA_WID*i) +: DATA_WID];
		end
	endgenerate
	
	//  -------------------------------------------------------------------------------------
	//	��Ϣ������M����
	//  -------------------------------------------------------------------------------------
	generate
		for(i=0; i<WORD_NUM; i=i+1) begin : m_data_word_reg_loop
			
			//	ģ������Ϊ0~15ʱ
			if(MODULE_INDEX < 16) begin
				
				//	��Ϣ��M���㹫ʽΪ M'(i) = M(i)��iȡֵ0~15
				always @ (posedge clk) begin
					
					//	��������Ϣ������M��Чʱ������
					if(i_m_data_vld) begin
						m_data_word_reg[i] <= m_data_word[i];
					end
				end
			end
			
			//	ģ������Ϊ16~63ʱ
			else begin
				
				//	��Ϣ����㹫ʽΪ M'(i) = M(i+1)��iȡֵ0~14
				if(i < 15) begin
					always @ (posedge clk) begin
					
						//	��������Ϣ������M��Чʱ������
						if(i_m_data_vld) begin
							m_data_word_reg[i] <= m_data_word[i+1];
						end
					end
				end
				
				//	��Ϣ����㹫ʽΪ M'(i) = rou1(M(i-1)) + M(i-6) + rou0(M(i-14)) + M(i-15)��iȡֵ15
				else begin
					always @ (posedge clk) begin
						
						//	��������Ϣ������M��Чʱ������
						if(i_m_data_vld) begin
							m_data_word_reg[i] <= rou1(m_data_word[i-1]) + m_data_word[i-6] + rou0(m_data_word[i-14]) + m_data_word[i-15];
						end
					end
				end
			end
		end
	endgenerate
	
	//  -------------------------------------------------------------------------------------
	//	�����Ϣ������Mƴ��
	//	����������Ϣ��M����32bit��wordΪ��λ������ƴ��
	//  -------------------------------------------------------------------------------------	
	generate
		for(i=0; i<WORD_NUM; i=i+1) begin : ov_m_data_loop
			assign	ov_m_data[(DATA_WID*i) +: DATA_WID] = m_data_word_reg[i];
		end
	endgenerate
	
	//  -------------------------------------------------------------------------------------
	//	�����չ��Ϣ������W
	//  -------------------------------------------------------------------------------------	
	generate
		//	ģ������Ϊ0~15ʱ
		if(MODULE_INDEX < 16) begin
			
			//	��չ��Ϣ��WΪ W = M(MODULE_INDEX)
			assign	ov_w_data = m_data_word_reg[MODULE_INDEX];
		end
		
		//	ģ������Ϊ16~63ʱ
		else begin
			
			//	��չ��Ϣ��WΪ W = M(15)
			assign	ov_w_data = m_data_word_reg[15];
		end
	endgenerate
	
	//  -------------------------------------------------------------------------------------
	//	�����Ϣ������M��Ч�������չ��Ϣ������W��Ч
	//  -------------------------------------------------------------------------------------	
	always @ (posedge clk) begin
		
		//	��λ
		if(rst) begin
			data_vld_reg <= 1'b0;
		end
		
		//	��������Ϣ������M��Ч����1��
		else begin
			data_vld_reg <= i_m_data_vld;
		end
	end
	
	assign o_m_data_vld = data_vld_reg;
	assign o_w_data_vld = data_vld_reg;
	
endmodule