//	********************************************************************************
//	ģ������clk_rst
//	��  �ܣ��������������ʱ�Ӻ͸�λ�ź�
//	��	Դ��
//	********************************************************************************
module clk_rst (
	
	//	�����ź�                                     	
	input	i_clk		,	//	����ʱ��

	//	����ź�
	output	o_clk		,	//	���ʱ��
	output	o_rst_sync		//	o_clkʱ���򣬸�λͬ��
	);
	
	
	//  ===============================================================================================
	//	�������źš�����˵��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�ź�˵��
	//  -------------------------------------------------------------------------------------
	wire	mmcm_locked	;	//	MMCM��ס	
		
		
	//  ===============================================================================================
	//	ʱ�ӡ���λģ������
	//  ===============================================================================================	
	//  -------------------------------------------------------------------------------------
	//	ʱ��ģ������
	//  -------------------------------------------------------------------------------------
	clk_gen clk_gen_inst(
		.i_clk			(i_clk			),	//	����ʱ��
		.o_clk			(o_clk			),	//	���ʱ��
		.o_mmcm_locked	(mmcm_locked	)	//	���MMCM����
	);
	
	//  -------------------------------------------------------------------------------------
	//	��λģ������
	//  -------------------------------------------------------------------------------------
	rst_sync rst_sync_inst(
		.clk				(o_clk			),	//	ģ�鹤��ʱ���ź�
		.i_rst_async		(~mmcm_locked	),	//	��λ�첽
		.i_rst_sync_en		(1'b1			),	//	��λͬ��ʹ��
		.o_rst_sync			(o_rst_sync		)	//	clkʱ���򣬸�λͬ��
	);
	
endmodule