//	********************************************************************************
//	ģ������uart_tx
//	��  �ܣ����ƴ��ڷ���
//	��	Դ��
//	********************************************************************************
module uart_tx # (
	
	//	�������
	parameter		IS_SIM			= "TRUE"		,	//	�Ƿ�Ϊ������ԣ�"TRUE" "FALSE"
	parameter		BAUD_RATE		= "115200"		,	//	�����ʣ�"9600" "115200"
	parameter		UART_DATA_WID	= 8					//	��������λ��8
	)                                                       	
	(                                                       	
	                                                        	
	//	ʱ�Ӹ�λ�ź�                                        	
	input							clk				,	//	ģ�鹤��ʱ���ź�
	input							rst				,	//	clkʱ���򣬸�λ
	                                                	
	//	�����ź�                                    	
	input	[UART_DATA_WID	-1:0]	iv_tx_data		,	//	clkʱ���򣬴��ڷ�������
	input							i_tx_data_vld	,	//	clkʱ���򣬴��ڷ���������Ч
	output							o_tx			,	//	clkʱ���򣬴��ڷ�����
	output							o_tx_done			//	clkʱ���򣬴��ڷ������
	);
	
	
	//  ===============================================================================================
	//	�������źš�����˵��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
	//	-----------------------------------------------------------------
	//	������λ��
	//	����16��λ����4��log2(16)=4
	//	-----------------------------------------------------------------
	function integer log2;
		
		//	�����ź�
		input	integer	data;
		
		//	�������� 
		integer data_tmp;
		
		//	�������  
		begin
			data_tmp = data - 1;
			for (log2=0; data_tmp>0; log2=log2+1) begin
				data_tmp = data_tmp >> 1;
			end
		end
	endfunction
	
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
	//	//	175MHz
//	localparam	BAUD_RATE_CNT_NUM	= (IS_SIM	 == "TRUE"	) ? 10		:
//									  (BAUD_RATE == "115200") ? 1519	: 
//									  (BAUD_RATE == "9600"  ) ? 18229	: 18229	;	//	�����ʼ�������������
	
	//	100MHz
	localparam	BAUD_RATE_CNT_NUM	= (IS_SIM	 == "TRUE"	) ? 10		:
									  (BAUD_RATE == "115200") ? 868		: 
									  (BAUD_RATE == "9600"  ) ? 10416	: 10416	;	//	�����ʼ�������������
	localparam	BAUD_RATE_CNT_WID	= log2(BAUD_RATE_CNT_NUM)					;	//	�����ʼ�����λ��
	localparam	BIT_CNT_NUM			= UART_DATA_WID + 2							;	//	bit��������������
	localparam	BIT_CNT_WID			= log2(BIT_CNT_NUM)							;	//	bit������λ��
	
	//  -------------------------------------------------------------------------------------
	//	�ź�˵��
	//  -------------------------------------------------------------------------------------
	//	�����ź�
	reg		[UART_DATA_WID		-1:0]	tx_data			= 'b0	;	//	clkʱ���򣬴��ڷ�������
	reg									tx_en			= 1'b0	;	//	clkʱ���򣬴��ڷ���ʹ��
	reg		[BAUD_RATE_CNT_WID	-1:0]	baud_rate_cnt	= 'b0	;	//	clkʱ���򣬲����ʼ�����
	reg		[BIT_CNT_WID		-1:0]	bit_cnt			= 'b0	;	//	clkʱ����bit������
	reg									tx						;	//	clkʱ���򣬴��ڷ�����
	
		
	//  ===============================================================================================
	//	���ڷ���
	//  ===============================================================================================	
	//  -------------------------------------------------------------------------------------
	//	���ڷ�����������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	�ڴ��ڷ���������Чʱ�����淢������
		if(i_tx_data_vld == 1'b1) begin
			tx_data <= iv_tx_data;
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	���ڷ���ʹ��
	//	��ʹFPGA��λ��ҲӦ�������������͸�PC���Է�ֹPC����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	�ڴ��ڷ���������Чʱ������ʹ��
		if(i_tx_data_vld == 1'b1) begin
			tx_en <= 1'b1;
		end
		
		//	�ڴ��ڷ������ʱ���õ�
		else if((tx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1))) begin
			tx_en <= 1'b0;
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	���ڲ����ʼ�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����ʹ����Чʱ������
		if(tx_en == 1'b1) begin
			
			//	�Ƶ����ֵ������
			if(baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) begin
				baud_rate_cnt <= 'b0;
			end
			
			//	�����ۼ�һ
			else begin
				baud_rate_cnt <= baud_rate_cnt + 1'b1;
			end
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	bit������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����ʹ����Ч���Ҳ����ʼ������Ƶ����ֵʱ������
		if((tx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1))) begin
			
			//	�Ƶ����ֵ������
			if(bit_cnt == (BIT_CNT_NUM - 1'b1)) begin
				bit_cnt <= 'b0;
			end
			
			//	�����ۼ�һ
			else begin
				bit_cnt <= bit_cnt + 1'b1;
			end
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	���ڷ�����
	//	��ʼλ0 + LSB + MSB + ֹͣλ1
	//  -------------------------------------------------------------------------------------
	always @ ( * ) begin
		
		//	�����ڼ�
		if(tx_en == 1'b1) begin
			
			//	����bit_cnt��ѡ��tx_data��Ӧ��bit����
			case(bit_cnt)
					
				//	��ʼλ0
				'd0	: begin
					tx = 1'b0;
				end
				
				//	tx_data��bit0-7
				'd1	,
				'd2	,
				'd3	,
				'd4	,
				'd5	,
				'd6	,
				'd7	,
				'd8	: begin
					tx = tx_data[bit_cnt-1'b1];
				end
				
				//	ֹͣλ1
				'd9	: begin
					tx = 1'b1;
				end
				
				//	����״̬����Ϊ1
				default	: begin
					tx = 1'b1;
				end
			endcase
		end
		
		//	�Ƿ����ڼ䣬���ָ�
		else begin
			tx = 1'b1;
		end
	end
	
	assign o_tx = tx;
	
	//  -------------------------------------------------------------------------------------
	//	���ڷ������
	//	����ʹ����Ч����bit�������Ƶ����ֵʱ���ø�
	//  -------------------------------------------------------------------------------------
	assign o_tx_done = ((tx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1))) ? 1'b1 : 1'b0;	
	
endmodule