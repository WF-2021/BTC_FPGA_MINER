//	********************************************************************************
//	ģ������rst_sync
//	��  �ܣ��첽��λͬ���ͷ�
//	��	Դ��
//	********************************************************************************
module rst_sync (
	
	//	�����ź�                                     	
	input	clk				,	//	ģ�鹤��ʱ���ź�
	input	i_rst_async		,	//	��λ�첽
	input	i_rst_sync_en	,	//	��λͬ��ʹ��

	//	����ź�
	output	o_rst_sync			//	clkʱ���򣬸�λͬ��
	);
	
	
	//  ===============================================================================================
	//	�������źš�����˵��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
	localparam	INITIALIZATION = 2'b11	;	//	��λͬ���Ĵ�����ʼֵ
	
	//  -------------------------------------------------------------------------------------
	//	�ź�˵��
	//  -------------------------------------------------------------------------------------
	wire	rst_sync_0	;	//	clkʱ���򣬸�λͬ��0
	wire	rst_sync_1	;	//	clkʱ���򣬸�λͬ��1
		
		
	//  ===============================================================================================
	//	�첽��λͬ���ͷ�
	//  ===============================================================================================	
	//  -------------------------------------------------------------------------------------
	//	FDPE�첽��λ�Ĵ���0
	//  -------------------------------------------------------------------------------------
	FDPE # (
		.INIT	(INITIALIZATION[0]	)	//	FDPE�����ʼֵ
	)
	fdpe_inst0 (
		.CE		(i_rst_sync_en		),	//	ʱ��ʹ��
		.C		(clk				),  //	ʱ��
		.PRE	(i_rst_async		),	//	�첽��λ����
		.D		(1'b0				),  //	�����ź�
		.Q		(rst_sync_0			)   //	����ź�
	);
	
	//  -------------------------------------------------------------------------------------
	//	FDPE�첽��λ�Ĵ���0
	//  -------------------------------------------------------------------------------------
	FDPE # (
		.INIT	(INITIALIZATION[1]	)	//	FDPE�����ʼֵ
	)
	fdpe_inst1 (
		.CE		(i_rst_sync_en		),	//	ʱ��ʹ��     
		.C		(clk				),	//	ʱ��         
		.PRE	(i_rst_async		),	//	�첽��λ���� 
		.D		(rst_sync_0			),	//	�����ź�     
		.Q		(rst_sync_1			) 	//	����ź�     
	);
	
	//  -------------------------------------------------------------------------------------
	//	��λͬ�����
	//  -------------------------------------------------------------------------------------
	assign o_rst_sync = rst_sync_1;
	
endmodule