//	********************************************************************************
//	ģ������uart_rx
//	��  �ܣ����ƴ��ڽ���
//	��	Դ��
//	********************************************************************************
module uart_rx # (
	
	//	�������
	parameter	IS_SIM				= "TRUE"		,	//	�Ƿ�Ϊ������ԣ�"TRUE" "FALSE"
	parameter	BAUD_RATE			= "115200"		,	//	�����ʣ�"9600" "115200"
	parameter	UART_DATA_WID		= 8				,	//	��������λ��8
	parameter	UART_RX_DATA_NUM	= 82				//	���ڽ��������ܸ�����82
	)                                                       	
	(                                                       	
	                                                        	
	//	ʱ�Ӹ�λ�ź�                                        	
	input							clk				,	//	ģ�鹤��ʱ���ź�
	input							rst				,	//	clkʱ���򣬸�λ

	//	�����ź�     
	input							i_rx			,	//	�첽ʱ���򣬴��ڽ�����
	output	[UART_DATA_WID	-1:0]	ov_rx_data		,	//	clkʱ���򣬴��ڽ�������
	output							o_rx_data_vld	,	//	clkʱ���򣬴��ڽ���������Ч	
	output							o_rx_busy			//	clkʱ���򣬴��ڽ���æµ
	);
	
	
	//  ===============================================================================================
	//	�������źš�����˵��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
	//	-----------------------------------------------------------------
	//	������λ��
	//	����16��λ����4��log2(16)=4
	//	-----------------------------------------------------------------
	function integer log2;
		
		//	�����ź�
		input	integer	data;
		
		//	�������� 
		integer data_tmp;
		
		//	�������  
		begin
			data_tmp = data - 1;
			for (log2=0; data_tmp>0; log2=log2+1) begin
				data_tmp = data_tmp >> 1;
			end
		end
	endfunction
	
	//  -------------------------------------------------------------------------------------
	//	����˵��
	//  -------------------------------------------------------------------------------------
//	//	175MHz
//	localparam	BAUD_RATE_CNT_NUM		= (IS_SIM	 == "TRUE"	) ? 10		:
//										  (BAUD_RATE == "115200") ? 1519	: 
//										  (BAUD_RATE == "9600"  ) ? 18229	: 18229	;	//	�����ʼ�������������
	
	//	100MHz
	localparam	BAUD_RATE_CNT_NUM		= (IS_SIM	 == "TRUE"	) ? 10		:
										  (BAUD_RATE == "115200") ? 868		: 
										  (BAUD_RATE == "9600"  ) ? 10416	: 10416	;	//	�����ʼ�������������
	localparam	BAUD_RATE_CNT_WID		= log2(BAUD_RATE_CNT_NUM)					;	//	�����ʼ�����λ��
	localparam	HALF_BAUD_RATE_CNT_NUM	= BAUD_RATE_CNT_NUM / 2						;	//	�벨���ʼ�������������
	localparam	BIT_CNT_NUM				= UART_DATA_WID + 2							;	//	bit��������������
	localparam	BIT_CNT_WID				= log2(BIT_CNT_NUM)							;	//	bit������λ��
	localparam	BYTE_CNT_NUM			= UART_RX_DATA_NUM							;	//	byte��������������
	localparam	BYTE_CNT_WID			= log2(BYTE_CNT_NUM)						;	//	byte������λ��
	
	//  -------------------------------------------------------------------------------------
	//	�ź�˵��
	//  -------------------------------------------------------------------------------------
	//	�����ź�	
	reg		[3					-1:0]	rx_dly			= 3'b111;	//	clkʱ���򣬴��ڽ����ߣ���1��	
	wire								rx_fall					;	//	clkʱ���򣬴��ڽ����ߣ��½���
	
	//	�����ź�
	reg									rx_en			= 1'b0	;	//	clkʱ���򣬴��ڽ���ʹ��
	reg		[BAUD_RATE_CNT_WID	-1:0]	baud_rate_cnt	= 'b0	;	//	clkʱ���򣬲����ʼ�����
	reg		[BIT_CNT_WID		-1:0]	bit_cnt			= 'b0	;	//	clkʱ����bit������
	reg		[BYTE_CNT_WID		-1:0]	byte_cnt		= 'b0	;	//	clkʱ����byte������
	reg		[UART_DATA_WID		-1:0]	rx_data			= 'b0	;	//	clkʱ���򣬴��ڽ�������
	reg									rx_busy			= 1'b0	;	//	clkʱ���򣬴��ڽ���æµ
	
		
	//  ===============================================================================================
	//	�����ź�
	//  ===============================================================================================	
	//  -------------------------------------------------------------------------------------
	//	�źŴ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		rx_dly <= {rx_dly, i_rx};
	end
	
	//  -------------------------------------------------------------------------------------
	//	�ź��������½���
	//  -------------------------------------------------------------------------------------
	assign rx_fall = ((rx_dly[1] == 1'b0) && (rx_dly[2] == 1'b1)) ? 1'b1 : 1'b0;
	
	
	//  ===============================================================================================
	//	���ڷ���
	//  ===============================================================================================	
	//  -------------------------------------------------------------------------------------
	//	���ڽ���ʹ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	���ڽ������½��أ�ʹ��
		if(rx_fall == 1'b1) begin
			rx_en <= 1'b1;
		end
		
		//	�ڴ��ڽ�����һ��byteʱ���õ�
		else if((rx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1))) begin
			rx_en <= 1'b0;
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	���ڲ����ʼ�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����ʹ����Чʱ������
		if(rx_en == 1'b1) begin
			
			//	�Ƶ����ֵ������
			if(baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) begin
				baud_rate_cnt <= 'b0;
			end
			
			//	�����ۼ�һ
			else begin
				baud_rate_cnt <= baud_rate_cnt + 1'b1;
			end
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	bit������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����ʹ����Ч���Ҳ����ʼ������Ƶ����ֵʱ������
		if((rx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1))) begin
			
			//	�Ƶ����ֵ������
			if(bit_cnt == (BIT_CNT_NUM - 1'b1)) begin
				bit_cnt <= 'b0;
			end
			
			//	�����ۼ�һ
			else begin
				bit_cnt <= bit_cnt + 1'b1;
			end
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	byte������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����ʹ����Ч����bit�������Ƶ����ֵʱ������
		if((rx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1))) begin
			
			//	�Ƶ����ֵ������
			if(byte_cnt == (BYTE_CNT_NUM - 1'b1)) begin
				byte_cnt <= 'b0;
			end
			
			//	�����ۼ�һ
			else begin
				byte_cnt <= byte_cnt + 1'b1;
			end
		end
	end
	
	//  -------------------------------------------------------------------------------------
	//	���ڽ�������
	//	��ʼλ0 + LSB + MSB + ֹͣλ1
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	����bit���������ڰ벨���ʴ����洮�ڽ�����
		if((rx_en == 1'b1) && (baud_rate_cnt == (HALF_BAUD_RATE_CNT_NUM - 1'b1)) && ((bit_cnt != 'b0) && (bit_cnt != (BIT_CNT_NUM - 1'b1)))) begin
			rx_data <= {i_rx, rx_data[UART_DATA_WID-1 : 1]};
		end
	end
	
	assign ov_rx_data = rx_data;
	
	//  -------------------------------------------------------------------------------------
	//	���ڽ���������Ч
	//	����ʹ����Ч����bit�������Ƶ����ֵʱ���ø�
	//  -------------------------------------------------------------------------------------
	assign o_rx_data_vld = ((rx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1))) ? 1'b1 : 1'b0;	
	
	//  -------------------------------------------------------------------------------------
	//	���ڽ���æµ
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		
		//	�ڴ��ڽ������½��ش����ø�
		if(rx_fall == 1'b1) begin
			rx_busy <= 1'b1;
		end
		
		//	����ʹ����Ч����byte�������Ƶ����ֵʱ���õ�
		else if((rx_en == 1'b1) && (baud_rate_cnt == (BAUD_RATE_CNT_NUM - 1'b1)) && (bit_cnt == (BIT_CNT_NUM - 1'b1)) && (byte_cnt == (BYTE_CNT_NUM - 1'b1))) begin
			rx_busy <= 1'b0;
		end
	end
	
	assign o_rx_busy = rx_busy;
	
endmodule